`include "utils.svh"

module system_tb();

  `TEST_PROGRAM test();

  test_harness `TH ();

endmodule
